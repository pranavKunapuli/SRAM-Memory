*** SPICE deck for cell basic_cell_read_write_stable{sch} from library memory
*** Created on Wed Nov 18, 2015 14:32:57
*** Last revised on Wed Nov 18, 2015 21:49:35
*** Written on Wed Nov 18, 2015 21:49:42 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include /home1/e/ese370/ptm/22nm_HP.pm

.global gnd vdd

*** TOP LEVEL CELL: basic_cell_read_write_stable{sch}
Mnmos@0 net@8 net@5 gnd gnd N L=0.022U W=0.022U
Mnmos@1 net@5 net@8 gnd gnd N L=0.022U W=0.022U
Mnmos@2 net@5 net@11 net@14 gnd N L=0.022U W=0.022U
Mnmos@3 net@20 net@11 net@8 gnd N L=0.022U W=0.022U
Mpmos@0 vdd net@5 net@8 vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@8 net@5 vdd P L=0.022U W=0.022U
VVPWL@0 net@14 gnd pwl (0ps 1v 110ps 1v 110ps 0v) DC 0V AC 0V 0
VVPWL@1 net@20 gnd pwl (0ps 0v 50ps 0v 50ps 1v) DC 0V AC 0V 0
VVPWL@2 net@11 gnd pwl (0ps 1v 10ps 1v 10ps 0v 50ps 0v 50ps 1v 100ps 1v 100ps 0v 110ps 0v 110ps 1v 120ps 1v 120ps 0v) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 1 AC 0
.END
