
.global gnd vdd

*** SUBCIRCUIT nor2 FROM CELL nor2{sch}
.SUBCKT nor2 A B O w=1
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O B gnd gnd N L=0.022U W=w*0.022U
Mnmos@1 O A gnd gnd N L=0.022U W=w*0.022U
Mpmos@0 vdd A net@23 vdd P L=0.022U W=w*2*0.022U
Mpmos@1 net@23 B O vdd P L=0.022U W=w*2*0.022U
.ENDS nor2

.END
