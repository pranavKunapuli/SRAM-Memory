
.include /home1/e/ese370/ptm/22nm_HP.pm
.include ./nand2.spi
.include ./nand3.spi

.global gnd vdd

*** SUBCIRCUIT full_tester FROM CELL full_tester{sch}
.SUBCKT full_tester full r0 r1 r2 r3 r4 r5 r6 r7 r8 w0 w1 w2 w3 w4 w5 w6 w7 w8
Xnand2@4 r0 w8 net@120 nand2 
Xnand2@5 r1 w0 net@124 nand2
Xnand2@6 r2 w1 net@122 nand2
Xnand2@7 r3 w2 net@128 nand2
Xnand2@14 r4 w3 net@126 nand2
Xnand2@9 r5 w4 net@130 nand2
Xnand2@15 r6 w5 net@131 nand2
Xnand2@11 r7 w6 net@132 nand2
Xnand2@13 r8 w7 net@136 nand2


Xnand3@0 net@120 net@124 net@122 net@140 nand3 w=2
Xnand3@1 net@128 net@126 net@130 net@138 nand3 w=2
Xnand3@2 net@131 net@132 net@136 net@142 nand3 w=2

Xnot@0 net@140 net@140n not w=4
Xnot@1 net@138 net@138n not w=4
Xnot@2 net@142 net@142n not w=4

Xnand3@3 net@140n net@138n net@142n full nand3 w=8
.ENDS full_tester

.END
