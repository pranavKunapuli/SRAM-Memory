
.global gnd vdd_clocking_clocking

*** SUBCIRCUIT not FROM CELL not{sch}
.SUBCKT not_clock A A_ w=1
** GLOBAL gnd
** GLOBAL vdd_clocking
Mnmos@0 A_ A gnd gnd N L=0.022U W=w*0.022U
Mpmos@0 vdd_clocking A A_ vdd_clocking P L=0.022U W=w*0.022U
.ENDS not

.END
