*** SPICE deck for cell sense_amp_test{sch} from library memory
*** Created on Wed Nov 18, 2015 23:16:08
*** Last revised on Wed Nov 18, 2015 23:57:17
*** Written on Wed Nov 18, 2015 23:59:09 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include /home1/e/ese370/ptm/22nm_HP.pm

*** SUBCIRCUIT memory__sense_amp FROM CELL sense_amp{sch}
.SUBCKT memory__sense_amp bit bit_b clk sense sense_b
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 sense_b sense net@25 gnd N L=0.022U W=0.044U
Mnmos@1 sense sense_b net@25 gnd N L=0.022U W=0.044U
Mnmos@4 net@25 clk gnd gnd N L=0.022U W=0.044U
Mpmos@0 bit clk sense vdd P L=0.022U W=0.088U
Mpmos@1 bit_b clk sense_b vdd P L=0.022U W=0.088U
Mpmos@2 vdd sense sense_b vdd P L=0.022U W=0.022U
Mpmos@3 vdd sense_b sense vdd P L=0.022U W=0.022U
.ENDS memory__sense_amp

.global gnd vdd

*** TOP LEVEL CELL: sense_amp_test{sch}
Mnmos@0 nmos@0_d net@29 nmos@0_s gnd N L=0.022U W=0.022U
Mnmos@1 nmos@1_d net@30 nmos@1_s gnd N L=0.022U W=0.022U
VVPWL@0 net@2 gnd pwl (0ps 0v 10ps 0v 10ps 1v 20ps 1v 20ps 0v 40ps 0v 40ps 1v) DC 0V AC 0V 0
VVPWL@1 net@9 gnd pwl (0ps 0.40v 30ps 0.40v 30ps 0.6v) DC 0V AC 0V 0
VVPWL@2 net@6 gnd pwl (0ps 0.6v 30ps 0.6v 30ps 0.40v) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 1 AC 0
Xsense_am@0 net@9 net@6 net@2 net@29 net@30 memory__sense_amp
.END
