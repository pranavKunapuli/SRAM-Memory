*** SPICE deck for cell v_ref_test{sch} from library memory
*** Created on Wed Nov 18, 2015 22:27:55
*** Last revised on Wed Nov 18, 2015 22:31:54
*** Written on Wed Nov 18, 2015 22:31:59 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include /home1/e/ese370/ptm/22nm_HP.pm

*** SUBCIRCUIT memory__v_ref FROM CELL v_ref{sch}
.SUBCKT memory__v_ref en out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@1 net@1 gnd gnd N L=0.022U W=0.088U
Mnmos@1 net@30 net@1 gnd gnd N L=0.022U W=0.352U
Mnmos@2 out en net@30 gnd N L=0.022U W=0.352U
Mpmos@0 vdd net@1 net@1 vdd P L=0.022U W=0.088U
Mpmos@1 vdd net@1 net@30 vdd P L=0.022U W=0.352U
.ENDS memory__v_ref

.global gnd vdd

*** TOP LEVEL CELL: v_ref_test{sch}
Rres@0 gnd net@5 1MEG
VVPWL@0 net@2 gnd pwl (0ps 0v 10ps 0v 10ps 1v 20ps 1v 20ps 0v 50ps 0v 50ps 1v) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 1 AC 0
Xv_ref@0 net@2 net@5 memory__v_ref
.END
