
.include ./column_precharger.spi
.include ./not_mem.spi

.global gnd vdd_mem

*** SUBCIRCUIT bit_driver FROM CELL bit_driver{sch}
.SUBCKT bit_driver bit bit_n in out precharge_en write_read_n

Mnmos@2 out_n out net@35 gnd N L=0.022U W=0.044U
Mnmos@3 out out_n net@35 gnd N L=0.022U W=0.044U
Mnmos@4 net@35 write_read_n gnd gnd N L=0.022U W=0.044U

Mnmos@5 bit write_read_n in gnd N L=0.022U W=0.352U
Mpmos@6 bit write_read_n out vdd_mem P L=0.022U W=0.022U

Mnmos@6 bit_n write_read_n in_n gnd N L=0.022U W=0.352U
Mpmos@7 bit_n write_read_n out_n vdd_mem P L=0.022U W=0.022U

Mpmos@4 vdd_mem out out_n vdd_mem P L=0.022U W=0.022U
Mpmos@5 vdd_mem out_n out vdd_mem P L=0.022U W=0.022U

Xcolumn_p@0 bit bit_n precharge_en column_precharger
Xnot_mem@0 in in_n not_mem
.ENDS bit_driver


.END
