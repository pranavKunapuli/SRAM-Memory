*** SPICE deck for cell basic_cell_read_write_tristate{sch} from library memory
*** Created on Wed Nov 18, 2015 13:34:12
*** Last revised on Thu Nov 19, 2015 10:54:54
*** Written on Thu Nov 19, 2015 10:55:04 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include /home1/e/ese370/ptm/22nm_HP.pm

*** SUBCIRCUIT memory__not FROM CELL not{sch}
.SUBCKT memory__not A A_ w=1
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 A_ A gnd gnd N L=0.022U W=w*0.022U
Mpmos@0 vdd A A_ vdd P L=0.022U W=w*0.022U
.ENDS memory__not

*** SUBCIRCUIT memory__sense_amp FROM CELL sense_amp{sch}
.SUBCKT memory__sense_amp bit bit_b clk sense sense_b
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 sense_b sense net@25 gnd N L=0.022U W=0.044U
Mnmos@1 sense sense_b net@25 gnd N L=0.022U W=0.044U
Mnmos@4 net@25 clk gnd gnd N L=0.022U W=0.044U
Mpmos@0 bit clk sense vdd P L=0.022U W=0.088U
Mpmos@1 bit_b clk sense_b vdd P L=0.022U W=0.088U
Mpmos@2 vdd sense sense_b vdd P L=0.022U W=0.022U
Mpmos@3 vdd sense_b sense vdd P L=0.022U W=0.022U
.ENDS memory__sense_amp

*** SUBCIRCUIT memory__sram FROM CELL sram{sch}
.SUBCKT memory__sram bit bit_b word
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@5 net@1 gnd gnd N L=0.022U W=0.022U
Mnmos@1 net@1 net@5 gnd gnd N L=0.022U W=0.022U
Mnmos@2 net@1 word bit gnd N L=0.022U W=0.022U
Mnmos@3 bit_b word net@5 gnd N L=0.022U W=0.022U
Mpmos@0 vdd net@1 net@5 vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@5 net@1 vdd P L=0.022U W=0.022U
.ENDS memory__sram

*** SUBCIRCUIT memory__tri_buffer FROM CELL tri_buffer{sch}
.SUBCKT memory__tri_buffer en in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out en net@5 gnd N L=0.022U W=0.352U
Mnmos@1 net@5 in gnd gnd N L=0.022U W=0.352U
Mpmos@0 net@4 net@1 out vdd P L=0.022U W=0.352U
Mpmos@1 vdd in net@4 vdd P L=0.022U W=0.352U
Xnot@0 en net@1 memory__not w=4
.ENDS memory__tri_buffer

*** SUBCIRCUIT memory__v_ref FROM CELL v_ref{sch}
.SUBCKT memory__v_ref out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@1 net@1 gnd gnd N L=0.022U W=0.088U
Mnmos@1 out net@1 gnd gnd N L=0.022U W=0.352U
Mpmos@0 vdd net@1 net@1 vdd P L=0.022U W=0.088U
Mpmos@1 vdd net@1 out vdd P L=0.022U W=0.352U
.ENDS memory__v_ref

.global gnd vdd

*** TOP LEVEL CELL: basic_cell_read_write_tristate{sch}
Mpmos@0 net@101 net@77 net@12 vdd P L=0.022U W=0.352U
Mpmos@1 net@101 net@77 net@7 vdd P L=0.022U W=0.352U
Mpmos@2 net@12 net@77 net@7 vdd P L=0.022U W=0.352U
VVPWL@0 net@0 gnd pwl (0ps 1v 20ps 1v 20ps 0v 40ps 0v 40ps 1v 80ps 1v 80ps 0v 100ps 0v 100ps 1v) DC 0V AC 0V 0
VVPWL@3 net@20 gnd pwl (0ps 1v 20ps 1v 20ps 0v 60ps 0v 60ps 1v 80ps 1v 80ps 0v) DC 0V AC 0V 0
VVPWL@4 net@77 gnd pwl (0ps 1v 20ps 1v 20ps 0v 40ps 0v 40ps 1v 80ps 1v 80ps 0v 100ps 0v 100ps 1v) DC 0V AC 0V 0
VVPWL@5 net@63 gnd pwl (0ps 1v 60ps 1v 60ps 0v) DC 0V AC 0V 0
VVPWL@6 net@147 gnd pwl (0v 1v 20ps 1v 20ps 0v 50ps 0v 50ps 1v 80ps 1v 80ps 0v 110ps 0v 110ps 1v) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 1 AC 0
Xnot@0 net@63 net@67 memory__not w=8
Xnot@2 net@152 not@2_A_ memory__not
Xnot@3 net@154 not@3_A_ memory__not
Xsense_am@0 net@7 net@12 net@147 net@152 net@154 memory__sense_amp
Xsram@0 net@7 net@12 net@0 memory__sram
Xtri_buff@0 net@20 net@63 net@7 memory__tri_buffer
Xtri_buff@1 net@20 net@67 net@12 memory__tri_buffer
Xv_ref@1 net@101 memory__v_ref
.END
