
.include /home1/e/ese370/ptm/22nm_HP.pm

.global gnd vdd

*** SUBCIRCUIT sense_amp FROM CELL sense_amp{sch}
.SUBCKT sense_amp bit bit_b clk sense sense_b w=1
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 sense_b sense s_gnd gnd N L=0.022U W=0.044U
Mnmos@1 sense sense_b s_gnd gnd N L=0.022U W=0.044U
Mnmos@4 s_gnd clk gnd gnd N L=0.022U W=0.044U
Mpmos@0 bit clk sense vdd P L=0.022U W=w*0.022U
Mpmos@1 bit_b clk sense_b vdd P L=0.022U W=w*0.022U
Mpmos@2 vdd sense sense_b vdd P L=0.022U W=0.022U
Mpmos@3 vdd sense_b sense vdd P L=0.022U W=0.022U
.ENDS sense_amp

.END
