
*** SUBCIRCUIT memory__not FROM CELL not{sch}
.SUBCKT memory__not A A_
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 A_ A gnd gnd N L=0.022U W=0.088U
Mpmos@0 vdd A A_ vdd P L=0.022U W=0.088U
.ENDS memory__not

.global gnd vdd

*** SUBCIRCUIT tri_buffer FROM CELL tri_buffer{sch}
.SUBCKT tri_buffer en in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out en net@5 gnd N L=0.022U W=0.352U
Mnmos@1 net@5 in gnd gnd N L=0.022U W=0.352U
Mpmos@0 net@4 net@1 out vdd P L=0.022U W=0.352U
Mpmos@1 vdd in net@4 vdd P L=0.022U W=0.352U
Xnot@0 en net@1 memory__not
.ENDS tri_buffer


Xtri_buffer en in out tri_buffer

.END
