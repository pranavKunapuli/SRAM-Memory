
.include /home1/e/ese370/ptm/22nm_HP.pm

.global gnd vdd_mem
.SUBCKT column_precharger bit bit_b en w=4

Mnmos@0 v_i v_i gnd gnd N L=0.022U W=w*0.25*0.022U
Mnmos@1 v_half v_i gnd gnd N L=0.022U W=w*0.022U
Mnmos@2 bit en v_half gnd N L=0.022U W=w*0.022U
Mnmos@3 bit_b en v_half gnd N L=0.022U W=w*0.022U
Mnmos@4 bit_b en bit gnd N L=0.022U W=w*0.022U
Mpmos@7 vdd_mem v_i v_i vdd_mem P L=0.022U W=w*0.25*0.022U
Mpmos@9 vdd_mem v_i v_half vdd_mem P L=0.022U W=w*0.022U
.ENDS column_precharger

.END
