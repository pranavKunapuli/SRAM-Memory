
.include /home1/e/ese370/ptm/22nm_HP.pm
.include ../bit_driver.spi
.include ../memory_column.spi
.include ../clock_delay.spi
.include ../not.spi
.include ../word_driver.spi
.include ../d_ff_sr.spi

.global gnd vdd

** GLOBAL gnd
** GLOBAL vdd
VVPWL@0 reset gnd pwl (0ns 1v 0ns 0v 1ns 0v 1ns 1v) DC 0V AC 0V 0
VVPWL@1 deq gnd pwl (0ns 0v 3.5ns 0v 3.5ns 1v) DC 0V AC 0V 0
VVPWL@2 enq gnd pwl (0ns 0v 1.5ns 0v 1.5ns 1v) DC 0V AC 0V 0
VVPWL@3 in gnd pwl (0ns 0v 3.8ns 0v 3.8ns 1v 5.8ns 1v 5.8ns 0v 7.8ns 0v 7.8ns 1v) DC 0V AC 0V 0
VVPulse@0 clk gnd pulse (0 1V 0ns 0ps 0ps 1ns 2ns) DC 0V AC 0V 0

VV_Generi@0 vdd gnd DC 1 AC 0
Xbit_driv@0 bit bit_b in_store out_store clk write_read_n bit_driver
Xclock_de@0 clk read_write_n clock_delay
Xmemory_c@0 bit bit_b w0 w1 w2 w3 w4 w5 w6 w7 w8 memory_column
Xnot@0 clk en not
Xnot@1 read_write_n write_read_n not
Xnot@2 out not@1_A_ not

Xword_dri@0 clk deq en enq read_write_n reset w0 w1 w2 w3 w4 w5 w6 w7 w8 empty full word_driver 

xd_ff_sr@0 clk empty empty_store net@xd_ff0 vdd vdd d_ff_sr
xd_ff_sr@1 clk full full_store net@xd_ff1 vdd vdd d_ff_sr

xd_ff_sr@2 clk in in_store net@xd_ff2 vdd vdd d_ff_sr
xd_ff_sr@3 clk out_store out net@xd_ff3 vdd vdd d_ff_sr

.ic v(bit)=0
.ic v(bit_b)=1

.END

plot xmemory_c@0.xsram@0.bit_i xmemory_c@0.xsram@1.bit_i xmemory_c@0.xsram@2.bit_i xmemory_c@0.xsram@3.bit_i 