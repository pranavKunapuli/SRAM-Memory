
.include /home1/e/ese370/ptm/22nm_HP.pm

.global gnd vdd
.SUBCKT column_precharger bit bit_b en_i w=4

Mnmos@0 v_i v_i gnd gnd N L=0.022U W=w*0.25*0.022U
Mnmos@1 v_half v_i gnd gnd N L=0.022U W=w*0.022U
Mnmos@2 bit en_i v_half gnd N L=0.022U W=w*0.022U
Mnmos@3 bit_b en_i v_half gnd N L=0.022U W=w*0.022U
Mnmos@4 bit_b en_i bit gnd N L=0.022U W=w*0.022U
Mpmos@7 vdd v_i v_i vdd P L=0.022U W=w*0.25*0.022U
Mpmos@9 vdd v_i v_half vdd P L=0.022U W=w*0.022U
.ENDS column_precharger

.END
