
.include /home1/e/ese370/ptm/22nm_HP.pm
.include ./nand3.spi

.global gnd vdd

*** SUBCIRCUIT d_ff_sr FROM CELL d_ff_sr{sch}
.SUBCKT d_ff_sr Clk D Q Q_ R S
** GLOBAL gnd
** GLOBAL vdd
Xnand3@4 S net@10 Q_ Q nand3
Xnand3@5 Q net@25 R Q_ nand3
Xnand3@6 S net@20 net@10 net@15 nand3
Xnand3@7 net@15 Clk R net@10 nand3
Xnand3@8 net@10 Clk net@20 net@25 nand3
Xnand3@9 net@25 D R net@20 nand3
.ENDS d_ff_sr

.END
