.include /home1/e/ese370/ptm/22nm_HP.pm

.global gnd vdd

*** SUBCIRCUIT not FROM CELL not{sch}
.SUBCKT not A A_ w=1
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 A_ A gnd gnd N L=0.022U W=w*0.022U
Mpmos@0 vdd A A_ vdd P L=0.022U W=w*0.022U
.ENDS not

.END
