
.include ./not_clock.spi
.include ./nand2.spi

.global gnd vdd_clocking

*** SUBCIRCUIT clock_delay FROM CELL clock_delay{sch}
.SUBCKT clock_delay clk clk_d
** GLOBAL gnd
** GLOBAL vdd_clocking
Xnand2@0 clk_n clk_n_d clk_d nand2 w=16
Xnot_clock@0 clk clk_n not_clock w=4

Xnot_clock@1 clk net@1 not_clock w=1
Xnot_clock@2 net@1 net@2 not_clock w=1
Xnot_clock@3 net@2 net@3 not_clock w=8
Xnot_clock@4 net@3 net@4 not_clock w=1
Xnot_clock@5 net@4 net@5 not_clock w=8
Xnot_clock@6 net@5 net@6 not_clock w=1
Xnot_clock@7 net@6 net@7 not_clock w=8
Xnot_clock@8 net@7 net@8 not_clock w=1
Xnot_clock@9 net@8 net@9 not_clock w=8
Xnot_clock@10 net@9 net@10 not_clock w=1
Xnot_clock@11 net@10 net@11 not_clock w=8
Xnot_clock@12 net@11 net@12 not_clock w=1
Xnot_clock@13 net@12 net@13 not_clock w=8
Xnot_clock@14 net@13 net@14 not_clock w=1
Xnot_clock@15 net@14 net@15 not_clock w=8
Xnot_clock@16 net@15 net@16 not_clock w=1
Xnot_clock@17 net@16 net@17 not_clock w=8
Xnot_clock@18 net@17 net@18 not_clock w=1
Xnot_clock@19 net@18 net@19 not_clock w=8
Xnot_clock@20 net@19 net@20 not_clock w=1
Xnot_clock@21 net@20 clk_n_d not_clock w=4

.ENDS clock_delay

.END
